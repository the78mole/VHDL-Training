-------------------------------------------------------------------------------
-- Title      : Configuration
-- Project    : ADS-Praktikum
-------------------------------------------------------------------------------
-- File       : config.vhd
-- Author     : Daniel Glaser
-- Company    : LfTE, FAU Erlangen-N�rnberg
-- Created    : 2006-07-03
-- Last update: 2006-07-03
-- Platform   : 
-- Standard   : VHDL'87
-------------------------------------------------------------------------------
-- Description: This file configures especially peripherial settings, some
--              modules need for proper configuration
-------------------------------------------------------------------------------
-- Copyright (c) 2006 LfTE, FAU Erlangen-N�rnberg
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author          Description
-- 2006-07-03  1.0      sidaglas	Created
-------------------------------------------------------------------------------

