-------------------------------------------------------------------------------
-- Title      : Multiplexer
-- Project    : ADS-Praktikum - 01_Multiplexer
-------------------------------------------------------------------------------
-- File       : multiplexer.vhd
-- Author     : Daniel Glaser
-- Company    : Lehrstuhl f�r Technische Elektronik, Universit�t Erlangen
-- Created    : 2006-06-27
-- Last update: 2006-07-10
-- Platform   : 
-- Standard   : VHDL'87
-------------------------------------------------------------------------------
-- Description: This module defines an 8-bit multiplexer for digital audio data
-------------------------------------------------------------------------------
-- Copyright (c) 2006 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author          Description
-- 2006-06-27  1.0      sidaglas        Created
-- 2006-06-27                           Finished
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;



entity multiplexer is

  port (

-- WRITE_HERE

    sel_s1 : in std_logic;
    sel_s2 : in std_logic);

end;



architecture multiplexer_behavioral of multiplexer is
begin


-- WRITE_HERE


end multiplexer_behavioral;


