

entity multiplexer is

  port (

-- WRITE_HERE

    sel_s1 : in std_logic;
    sel_s2 : in std_logic);

end;


